// File: vga_example.sv
// This is the top level design for EE178 Lab #4.

// The `timescale directive specifies what the
// simulation time units are (1 ns here) and what
// the simulator time step should be (1 ps here).

`timescale 1 ns / 1 ps

// Declare the module and its ports.

module vga_example (
  input  logic clk,
  output logic vs,
  output logic hs,
  output logic [3:0] r,
  output logic [3:0] g,
  output logic [3:0] b,
  output logic pclk_mirror
  );

  // Converts 100 MHz clk into 40 MHz pclk.
  // This uses a vendor specific primitive
  // called MMCME2, for frequency synthesis.

  logic clk_in;
  logic locked;
  logic clk_fb;
  logic clk_ss;
  logic clk_out;
  logic pclk;
  (* KEEP = "TRUE" *) 
  (* ASYNC_REG = "TRUE" *)
  logic [7:0] safe_start = 0;

  IBUF clk_ibuf (.I(clk),.O(clk_in));

  MMCME2_BASE #(
    .CLKIN1_PERIOD(10.000),
    .CLKFBOUT_MULT_F(10.000),
    .CLKOUT0_DIVIDE_F(25.000))
  clk_in_mmcme2 (
    .CLKIN1(clk_in),
    .CLKOUT0(clk_out),
    .CLKOUT0B(),
    .CLKOUT1(),
    .CLKOUT1B(),
    .CLKOUT2(),
    .CLKOUT2B(),
    .CLKOUT3(),
    .CLKOUT3B(),
    .CLKOUT4(),
    .CLKOUT5(),
    .CLKOUT6(),
    .CLKFBOUT(clkfb),
    .CLKFBOUTB(),
    .CLKFBIN(clkfb),
    .LOCKED(locked),
    .PWRDWN(1'b0),
    .RST(1'b0)
  );

  BUFH clk_out_bufh (.I(clk_out),.O(clk_ss));
  always_ff @(posedge clk_ss) safe_start<= {safe_start[6:0],locked};

  BUFGCE clk_out_bufgce (.I(clk_out),.CE(safe_start[7]),.O(pclk));

  // Mirrors pclk on a pin for use by the testbench;
  // not functionally required for this design to work.

  ODDR pclk_oddr (
    .Q(pclk_mirror),
    .C(pclk),
    .CE(1'b1),
    .D1(1'b1),
    .D2(1'b0),
    .R(1'b0),
    .S(1'b0)
  );

  // Instantiate the vga_timing module, which is
  // the module you are designing for this lab.

  logic [10:0] vcount, hcount;
  logic vsync, hsync;
  logic vblnk, hblnk;

  vga_timing my_timing (
    .vcount(vcount),
    .vsync(vsync),
    .vblnk(vblnk),
    .hcount(hcount),
    .hsync(hsync),
    .hblnk(hblnk),
    .pclk(pclk)
  );

  // This is a simple test pattern generator.
  
  always_ff @(posedge pclk)
  begin
    // Just pass these through.
    hs <= hsync;
    vs <= vsync;
    // During blanking, make it it black.
    if (vblnk || hblnk) {r,g,b} <= 12'h0_0_0; 
    else
    begin
      // Active display, top edge, make a yellow line.
      if (vcount == 0) {r,g,b} <= 12'hf_f_0;
      // Active display, bottom edge, make a red line.
      else if (vcount == 599) {r,g,b} <= 12'hf_0_0;
      // Active display, left edge, make a green line.
      else if (hcount == 0) {r,g,b} <= 12'h0_f_0;
      // Active display, right edge, make a blue line.
      else if (hcount == 799) {r,g,b} <= 12'h0_0_f;
      // Active display, interior, fill with gray.
      // You will replace this with your own test.

      //my logo 
      else if((150<vcount)&&(vcount<250)&&(320<hcount)&&(hcount<330)) begin //N
        {r,g,b} <= 12'hf_f_0;
      end

      else if ((330<hcount)&&(hcount<390)&&(170<vcount)&&(vcount<180))begin //N
        {r,g,b} <= 12'hf_f_0;

      end
      else if ((390<hcount)&&(hcount<400)&&(170<vcount)&&(vcount<250))begin
        {r,g,b} <= 12'hf_f_0;
      end

      else if ((500<hcount)&&(hcount<510)&&(150<vcount)&&(vcount<250))begin
        {r,g,b} <= 12'hf_f_0;
      end
      else if((510<hcount)&&(hcount<570)&&(130<vcount)&&(vcount<140))begin
        {r,g,b} <= 12'hf_f_0;
      end
      // //skos
      // else if((510<=hcount<=570)&&(140<=vcount<=250))begin
      //   if((510<hcount<515)&&(140<vcount<150))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((515<=hcount<520)&&(150<=vcount<160))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((520<=hcount<525)&&(160<=vcount<170))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((525<=hcount<530)&&(170<=vcount<180))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((530<=hcount<535)&&(180<=vcount<190))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((535<=hcount<540)&&(190<=vcount<200))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((540<=hcount<545)&&(200<=vcount<210))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((545<=hcount<550)&&(210<=vcount<220))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((550<=hcount<555)&&(220<=vcount<230))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((555<=hcount<560)&&(230<=vcount<240))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else if((560<=hcount<570)&&(240<=vcount<250))begin
      //     {r,g,b} <= 12'hf_f_0;
      //   end
      //   else {r,g,b} <= 12'h8_8_8;  
      // end
      
      else {r,g,b} <= 12'h8_8_8;    
    end
  end

endmodule
